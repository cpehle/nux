module Syn_io_dummy
  ( input logic clk, reset,
    Syn_io_if.syn syn_io);


endmodule
